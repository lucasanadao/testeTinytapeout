/*
 * Copyright (c) 2024 Lucas Augusto dos Santos Anadão
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

// just a stub to keep the Tiny Tapeout tools happy

module tt_um_teste_tinytapeout (
    input  wire [7:0] ui_in,
    output wire [7:0] uo_out,
    input  wire [7:0] uio_in,
    output wire [7:0] uio_out,
    output wire [7:0] uio_oe,
    input  wire       ena,
    input  wire       clk,
    input  wire       rst_n
);

endmodule
